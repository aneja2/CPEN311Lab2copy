module tb_task2();

// Your testbench goes here. Our toplevel will give up after 1,000,000 ticks.

endmodule: tb_task2
